`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/27/2022 03:00:06 PM
// Design Name: 
// Module Name: HIDtest
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module HIDtest();
reg kbdclk;
reg kbddat;
reg clk;
wire [7:0] decoded;
wire [4:0] kbout;
wire state;
HID h(kbdclk,kbddat,decoded);
kbdWrapper k(clk,kbdclk,kbddat,kbout,state);
initial begin
//should transmit F0 followed by 2B (keycode F)
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
kbdclk=1;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=0;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
kbdclk=1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
kbddat=1;
kbdclk=0;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;
clk=1;
#1;
clk=0;
#1;


end
endmodule

